module char_rom(
  input        [6:0] addr,
  output reg [127:0] data_out
);


always @(*) begin
  case (addr)
  default: data_out = 128'hffffffffffffffffffffffffffffffff;
    8'h00: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h01: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h02: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h03: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h04: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h05: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h06: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h07: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h08: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h09: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h0A: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h0B: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h0C: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h0D: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h0E: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h0F: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h10: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h11: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h12: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h13: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h14: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h15: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h16: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h17: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h18: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h19: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h1A: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h1B: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h1C: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h1D: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h1E: data_out = 128'hffffffffffffffffffffffffffffffff;
	 8'h1F: data_out = 128'hffffffffffffffffffffffffffffffff;
    /* U+20 " " */
    8'h20: data_out = 128'h00000000000000000000000000000000;
	 /* U+21 "!" */
	 8'h21: data_out = 128'h00001010101010101000101000000000;
    /* U+22 "\"" */
    8'h22: data_out = 128'h00242424000000000000000000000000;
    /* U+23 "#" */
    8'h23: data_out = 128'h00002424247e24247e24242400000000;
    /* U+24 "$" */
    8'h24: data_out = 128'h0010107c9290907c1212927c10100000;
    /* U+25 "%" */
    8'h25: data_out = 128'h0000649468081010202c524c00000000;
    /* U+26 "&" */
    8'h26: data_out = 128'h000018242418304a4444443a00000000;
    /* U+27 "'" */
    8'h27: data_out = 128'h00101010000000000000000000000000;
    /* U+28 "(" */
    8'h28: data_out = 128'h00000810202020202020100800000000;
    /* U+29 ")" */
    8'h29: data_out = 128'h00002010080808080808102000000000;
    /* U+2A "*" */
    8'h2A: data_out = 128'h000000000024187e1824000000000000;
    /* U+2B "+" */
    8'h2B: data_out = 128'h000000000010107c1010000000000000;
    /* U+2C "," */
    8'h2C: data_out = 128'h00000000000000000000101020000000;
    /* U+2D "-" */
    8'h2D: data_out = 128'h000000000000007e0000000000000000;
    /* U+2E "." */
    8'h2E: data_out = 128'h00000000000000000000101000000000;
    /* U+2F "/" */
    8'h2F: data_out = 128'h00000404080810102020404000000000;
    /* U+30 "0" */
    8'h30: data_out = 128'h00003c4242464a526242423c00000000;
    /* U+31 "1" */
    8'h31: data_out = 128'h00000818280808080808083e00000000;
    /* U+32 "2" */
    8'h32: data_out = 128'h00003c42420204081020407e00000000;
    /* U+33 "3" */
    8'h33: data_out = 128'h00003c4242021c020242423c00000000;
    /* U+34 "4" */
    8'h34: data_out = 128'h000002060a1222427e02020200000000;
    /* U+35 "5" */
    8'h35: data_out = 128'h00007e4040407c020202423c00000000;
    /* U+36 "6" */
    8'h36: data_out = 128'h00001c2040407c424242423c00000000;
    /* U+37 "7" */
    8'h37: data_out = 128'h00007e02020404080810101000000000;
    /* U+38 "8" */
    8'h38: data_out = 128'h00003c4242423c424242423c00000000;
    /* U+39 "9" */
    8'h39: data_out = 128'h00003c424242423e0202043800000000;
    /* U+3A ":" */
    8'h3A: data_out = 128'h00000000001010000000101000000000;
    /* U+3B ";" */
    8'h3B: data_out = 128'h00000000001010000000101020000000;
    /* U+3C "<" */
    8'h3C: data_out = 128'h00000004081020402010080400000000;
    /* U+3D "=" */
    8'h3D: data_out = 128'h00000000007e00007e00000000000000;
    /* U+3E ">" */
    8'h3E: data_out = 128'h00000040201008040810204000000000;
    /* U+3F "?" */
    8'h3F: data_out = 128'h00003c42424204080800080800000000;
    /* U+40 "@" */
    8'h40: data_out = 128'h00007c829ea2a2a2a69a807e00000000;
    /* U+41 "A" */
    8'h41: data_out = 128'h00003c424242427e4242424200000000;
    /* U+42 "B" */
    8'h42: data_out = 128'h00007c4242427c424242427c00000000;
    /* U+43 "C" */
    8'h43: data_out = 128'h00003c42424040404042423c00000000;
    /* U+44 "D" */
    8'h44: data_out = 128'h00007844424242424242447800000000;
    /* U+45 "E" */
    8'h45: data_out = 128'h00007e40404078404040407e00000000;
    /* U+46 "F" */
    8'h46: data_out = 128'h00007e40404078404040404000000000;
    /* U+47 "G" */
    8'h47: data_out = 128'h00003c424240404e4242423c00000000;
    /* U+48 "H" */
    8'h48: data_out = 128'h0000424242427e424242424200000000;
    /* U+49 "I" */
    8'h49: data_out = 128'h00003810101010101010103800000000;
    /* U+4A "J" */
    8'h4A: data_out = 128'h00000e04040404040444443800000000;
    /* U+4B "K" */
    8'h4B: data_out = 128'h00004244485060605048444200000000;
    /* U+4C "L" */
    8'h4C: data_out = 128'h00004040404040404040407e00000000;
    /* U+4D "M" */
    8'h4D: data_out = 128'h000082c6aa9292828282828200000000;
    /* U+4E "N" */
    8'h4E: data_out = 128'h000042424262524a4642424200000000;
    /* U+4F "O" */
    8'h4F: data_out = 128'h00003c42424242424242423c00000000;
    /* U+50 "P" */
    8'h50: data_out = 128'h00007c424242427c4040404000000000;
    /* U+51 "Q" */
    8'h51: data_out = 128'h00003c424242424242424a3c02000000;
    /* U+52 "R" */
    8'h52: data_out = 128'h00007c424242427c5048444200000000;
    /* U+53 "S" */
    8'h53: data_out = 128'h00003c4240403c020242423c00000000;
    /* U+54 "T" */
    8'h54: data_out = 128'h0000fe10101010101010101000000000;
    /* U+55 "U" */
    8'h55: data_out = 128'h00004242424242424242423c00000000;
    /* U+56 "V" */
    8'h56: data_out = 128'h00004242424242242424181800000000;
    /* U+57 "W" */
    8'h57: data_out = 128'h000082828282829292aac68200000000;
    /* U+58 "X" */
    8'h58: data_out = 128'h00004242242418182424424200000000;
    /* U+59 "Y" */
    8'h59: data_out = 128'h00008282444428101010101000000000;
    /* U+5A "Z" */
    8'h5A: data_out = 128'h00007e02020408102040407e00000000;
    /* U+5B "[" */
    8'h5B: data_out = 128'h00003820202020202020203800000000;
    /* U+5C "\\" */
    8'h5C: data_out = 128'h00004040202010100808040400000000;
    /* U+5D "]" */
    8'h5D: data_out = 128'h00003808080808080808083800000000;
    /* U+5E "^" */
    8'h5E: data_out = 128'h00102844000000000000000000000000;
    /* U+5F "_" */
    8'h5F: data_out = 128'h000000000000000000000000007e0000;
    /* U+60 "`" */
    8'h60: data_out = 128'h10080000000000000000000000000000;
    /* U+61 "a" */
    8'h61: data_out = 128'h00000000003c023e4242423e00000000;
    /* U+62 "b" */
    8'h62: data_out = 128'h00004040407c42424242427c00000000;
    /* U+63 "c" */
    8'h63: data_out = 128'h00000000003c42404040423c00000000;
    /* U+64 "d" */
    8'h64: data_out = 128'h00000202023e42424242423e00000000;
    /* U+65 "e" */
    8'h65: data_out = 128'h00000000003c42427e40403c00000000;
    /* U+66 "f" */
    8'h66: data_out = 128'h00000e10107c10101010101000000000;
    /* U+67 "g" */
    8'h67: data_out = 128'h00000000003e42424242423e02023c00;
    /* U+68 "h" */
    8'h68: data_out = 128'h00004040407c42424242424200000000;
    /* U+69 "i" */
    8'h69: data_out = 128'h00001010003010101010103800000000;
    /* U+6A "j" */
    8'h6A: data_out = 128'h00000404000c04040404040444443800;
    /* U+6B "k" */
    8'h6B: data_out = 128'h00004040404244487048444200000000;
    /* U+6C "l" */
    8'h6C: data_out = 128'h00003010101010101010103800000000;
    /* U+6D "m" */
    8'h6D: data_out = 128'h0000000000fc92929292929200000000;
    /* U+6E "n" */
    8'h6E: data_out = 128'h00000000007c42424242424200000000;
    /* U+6F "o" */
    8'h6F: data_out = 128'h00000000003c42424242423c00000000;
    /* U+70 "p" */
    8'h70: data_out = 128'h00000000007c42424242427c40404000;
    /* U+71 "q" */
    8'h71: data_out = 128'h00000000003e42424242423e02020200;
    /* U+72 "r" */
    8'h72: data_out = 128'h00000000005e60404040404000000000;
    /* U+73 "s" */
    8'h73: data_out = 128'h00000000003e40403c02027c00000000;
    /* U+74 "t" */
    8'h74: data_out = 128'h00001010107c10101010100e00000000;
    /* U+75 "u" */
    8'h75: data_out = 128'h00000000004242424242423e00000000;
    /* U+76 "v" */
    8'h76: data_out = 128'h00000000004242422424181800000000;
    /* U+77 "w" */
    8'h77: data_out = 128'h00000000008282929292927c00000000;
    /* U+78 "x" */
    8'h78: data_out = 128'h00000000004242241824424200000000;
    /* U+79 "y" */
    8'h79: data_out = 128'h00000000004242424242423e02023c00;
    /* U+7A "z" */
    8'h7A: data_out = 128'h00000000007e04081020407e00000000;
    /* U+7B "{" */
    8'h7B: data_out = 128'h00000c10101020101010100c00000000;
    /* U+7C "|" */
    8'h7C: data_out = 128'h00001010101010101010101000000000;
    /* U+7D "}" */
    8'h7D: data_out = 128'h00003008080804080808083000000000;
    /* U+7E "~" */
    8'h7E: data_out = 128'h0062928c000000000000000000000000;
	 8'h7F: data_out = 128'hffffffffffffffffffffffffffffffff;
  endcase
end

endmodule